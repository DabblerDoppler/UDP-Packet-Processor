
const logic [3:0] IP_VERSION = 4;
//the desired header length is 20 or greater, but we multiply
//ip_header_length by 4, so it's really 5 or greater.
const logic [3:0] HEADER_LENGTH = 5;

module filter_core(
    //the filter's combinational, but the configuration module requires these.
    input logic clk, rst_n,
    // Header data input
    input logic [511:0] data,

    // AXI style configuration interface
    input  logic         cfg_we,
    input  logic  [3:0]  cfg_waddr,
    input  logic [31:0]  cfg_wdata,
    input  logic  [3:0]  cfg_raddr,
    output logic [31:0]  cfg_rdata,

    output logic filters_valid
);
    logic eth_valid, ip_valid, udp_valid;

    filter_config my_configuration (.clk, .rst_n, 
    .cfg_we, .cfg_waddr, .cfg_wdata, .cfg_raddr, .cfg_rdata, 
    .local_mac(cfg_local_mac), .ethertype(cfg_ethertype), 
    .ip_protocol(cfg_ip_protocol), .ip_base(cfg_ip_base), .ip_mask(cfg_ip_mask), 
    .udp_dst_port(cfg_dest_port));

    //Ethernet logic.
    logic [47:0] dest_mac, cfg_local_mac;
    logic [15:0] ethertype, cfg_ethertype;
    
    assign dest_mac = data[47:0];
    assign ethertype = data[111:96];

    assign eth_valid = (dest_mac == cfg_local_mac &&
            ethertype == cfg_ethertype);

    //IP logic - this contains most of our filtering.
    logic [3:0] ip_version, ip_header_length;
    logic [7:0] ip_protocol, cfg_ip_protocol;
    logic [31:0] ip_dest;

    assign ip_version = data[115:112];
    assign ip_header_length = data[119:116];
    assign ip_protocol = data[191:184];
    assign ip_dest = data[255:224];

    assign version_correct = ip_version == IP_VERSION;
    assign header_length_correct = ip_header_length == HEADER_LENGTH;
    assign protocol_correct = ip_protocol == cfg_ip_protocol;
    //bitwise AND the destination IP and our config mask, and compare that to the base.
    assign dest_correct = (ip_dest & cfg_ip_mask) == cfg_ip_base;

    assign ip_valid = (version_correct && 
                        header_length_correct && 
                        protocol_correct && 
                        dest_correct)

    //UDP logic
    logic [15:0] dest_port, cfg_dest_port;

    assign dest_port = data[388:303];

    assign udp_valid = (dest_port == cfg_dest_port);

    //Overall, the data is valid only if all our filters validate it.
    assign filters_valid = (eth_valid && ip_valid && udp_valid);
        
endmodule